`timescale 1ns/1ps
`default_nettype none

module :VIM_EVAL:expand("<afile>:t:r"):END_EVAL: (
);

endmodule

`resetall
