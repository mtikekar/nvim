module :VIM_EVAL:expand("<afile>:t:r"):END_EVAL: #() (
);

endmodule
